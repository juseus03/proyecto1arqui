//---------------------------------------------------------------------------
// SharkBoad ExampleModule
// Fredy Segura Q.
// Josnelihurt Rodriguez Barajas
// fsegura@uniandes.edu.co
// j.rodriguez52@uniandes.edu.co
// Top Level Design for the Xilinx Spartan 3-100E Device
//---------------------------------------------------------------------------

/*#
# SharkBoad
# Copyright (C) 2012 Bogotá, Colombia
#
# This program is free software: you can redistribute it and/or modify
# it under the terms of the GNU General Public License as published by
# the Free Software Foundation, version 3 of the License.
#
# This program is distributed in the hope that it will be useful,
# but WITHOUT ANY WARRANTY; without even the implied warranty of
# MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
# GNU General Public License for more details.
#
# You should have received a copy of the GNU General Public License
# along with this program.  If not, see <http://www.gnu.org/licenses/>.
#*/

module decoder #(
	parameter SELECTION = 4,		//NUMBER OF SELECTION BITS
	parameter DATAWIDTH = 9
	)
	(
	input			[SELECTION-1:0] 	sSelDeco,
	output reg		[DATAWIDTH-1:0] 	sOutDeco
	);
	always@(*)
	begin
	case (sSelDeco)	
		3'b000: sOutDeco = 8'b11111110;//R0
		3'b001: sOutDeco = 8'b11111101;//R1
		3'b010: sOutDeco = 8'b11111011;//R2
		3'b011: sOutDeco = 8'b11110111;//R3
		3'b100: sOutDeco = 8'b11101111;//R4
		3'b101: sOutDeco = 8'b11011111;//RP0
		3'b110: sOutDeco = 8'b10111111;//RP1
		3'b111: sOutDeco = 8'b11111111; //Not register selected to write
		default :   sOutDeco = 8'b1111110; //
		endcase
	end
endmodule
